--MICHAEL LOWE 
--EEL 4712 LAB 2 PART 2

library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all;
 



entity alu_ns is
	
	
	generic(
		
			WIDTH: positive := 16
	);
	
	
	
	port(
			input1: in std_logic_vector(WIDTH-1 downto 0); 
			input2: in std_logic_vector(WIDTH-1 downto 0);
			sel: in std_logic_vector(3 downto 0);
			output: out std_logic_vector(WIDTH-1 downto 0);
			overflow: out std_logic
	);	 
	
end alu_ns; 


architecture ALU of alu_ns is
	
	--Declare mux select lines as constants for the duration of process
	
	constant C_ADD: std_logic_vector(3 downto 0) := "0000";
	constant C_SUB: std_logic_vector(3 downto 0) := "0001"; 
	constant C_MULT: std_logic_vector(3 downto 0) := "0010"; 
	constant C_AND: std_logic_vector(3 downto 0) := "0011"; 
	constant C_OR: std_logic_vector(3 downto 0) := "0100"; 
	constant C_XOR: std_logic_vector(3 downto 0) := "0101"; 
	constant C_NOR: std_logic_vector(3 downto 0) := "0110"; 
	constant C_NOT: std_logic_vector(3 downto 0) := "0111"; 
	constant C_shift_left: std_logic_vector(3 downto 0) := "1000"; 
	constant C_shift_right: std_logic_vector(3 downto 0) := "1001"; 
	constant C_swap_bits: std_logic_vector(3 downto 0) := "1010";
	constant C_reverse_bits: std_logic_vector(3 downto 0) := "1011"; 
	constant C_whatever: std_logic_vector(3 downto 0) := "1111"; 
	
begin
	
	--BEGIN short circuit evaluation 
	process(sel, input1, input2)
		
		variable temp : unsigned(WIDTH-1 downto 0);
		variable operation_res : unsigned(2*WIDTH -1 downto 0) := (others=> '0');
		variable operation_res_2: unsigned(WIDTH downto 0) :=  (others => '0'); 
		 
			
	begin
		
		case sel is
			
		--ADDITION 		
		when C_ADD => 
			
			temp := unsigned(input1) + unsigned(input2);
			for i in 0 to (WIDTH -1 ) loop
			
				if(temp(i) = '1')
					then overflow <= '1';
				else
					overflow <= '0'; 
				end if; 
				
		end loop; 
			 
			
		--SUBTRACTION 
		when C_SUB =>
			
			temp := unsigned(input1) - unsigned(input2); 
			
			for i in  0 to (WIDTH-1) loop
			
				if(temp(i) = '1')
					then overflow <= '1'; 
				else
					overflow <= '0'; 
				end if; 
				
		end loop; 
			
			
		
		--MULTIPLICATION
				
	when C_MULT =>
		operation_res := unsigned(input1) * unsigned(input2);
		for i in (WIDTH -1) to (WIDTH*2 -1) loop
		
			if(operation_res(i) = '1')
				then overflow <= '1'; 
			else
					overflow <= '0'; 
			end if;
			 
		end loop; 
		
		temp := operation_res(WIDTH-1 downto 0); 
		
	when C_AND =>
		temp := unsigned((input1) AND (input2));
		overflow <= '0';  
		
	when C_OR =>
		temp := unsigned((input1) OR (input2)); 
		overflow <= '0';
		
	when C_XOR =>
		temp := unsigned((input1) XOR (input2));
		overflow <= '0';
		 
	when C_NOR =>
		temp := unsigned((input1) NOR (input2));
		overflow <= '0';
		 
	when C_NOT =>
		temp := unsigned( not ((input1)));
		overflow <= '0'; 

		
	when C_shift_left => 
		
		temp := SHIFT_LEFT(unsigned(input1), 1);
		
		if(input1(WIDTH-1) = '1')
			then overflow <= '1';
		else
		overflow <= '0';	
		end if;
		
		
	when C_shift_right =>
		temp := SHIFT_RIGHT(unsigned(input1), 1); 
		overflow <= '0';
		
		
	when C_swap_bits =>
		if(WIDTH mod 2 = 0)
			then temp := SHIFT_RIGHT(unsigned(input1), WIDTH/2) OR SHIFT_LEFT(unsigned(input2), WIDTH/2);
		else
			temp:= SHIFT_RIGHT(unsigned(input1), WIDTH/2 +1) OR SHIFT_LEFT(unsigned(input2), WIDTH/2 -1);
		end if; 
		overflow <= '0';
	
	
	--Iterates from vector of size length backwards and assigns to temp forwards. 
	when C_reverse_bits =>
		for i in 0 to WIDTH-1 loop
			temp(i) := input1((WIDTH-1) - i);
		end loop;

	when C_whatever =>

		operation_res_2 := unsigned((resize(not(unsigned(input1)), WIDTH +1))) + resize(unsigned(input2), WIDTH +1); 

			if(operation_res_2(WIDTH) = '1')
				then overflow <= '1'; 
			end if; 
				

		temp := operation_res_2(WIDTH-1 downto 0); 



		
	--TBA when other functions are needed  
	when others => null;
		
		--overflow <= '0';
		
		end case;
		
		
		
		output <= std_logic_vector(temp); 
		 

	end process; 
end ALU;

	